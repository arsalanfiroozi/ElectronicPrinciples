Lab4 - Arsalan Firoozi 97102225

***************** DC *************************
VCC 100 0 10
VEE 200 0 -10

***************** Resistors ******************
R2 1 0 455
R1 2 1 455
R3 2 3 455
C1 3 4 1u
Vinitial 4 0 5v

***************** Opamp **********************
Eopamp 2 0 1 3 MAX=10 MIN=-10 10000

.op
.tran 1n 18ms

.end